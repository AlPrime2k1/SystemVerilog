///////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Company: Scaledge Technology
// Engineer: Kirti Kumar
// 
// Module Name: fifo_defines
// Project Name: FIFO Verification
// Description: Definitions for fifo
///////////////////////////////////////////////////////////////////////////////////////////////////////////////

`ifndef FIFO_DEFINES_SV
`define FIFO_DEFINES_SV
`define PTR		   4

`define DATA_WIDTH 8
`define DEPTH 	   8
`define GAP		   2

`endif
