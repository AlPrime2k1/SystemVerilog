//////////////////////////////////////////////////////////////////////////////////
// Company: Scaledge Technology
// Engineer: Kirti Kumar
// 
// Module Name: ram_defines
// Project Name: RAM Verification
// Description: This file consists of definitions used throughout the project
//////////////////////////////////////////////////////////////////////////////////

`ifndef RAM_DEFINES_SV
`define RAM_DEFINES_SV

`define ADDR_WIDTH 4
`define DATA_WIDTH 8
`define DEPTH 	   16

`endif