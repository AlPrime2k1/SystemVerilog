library verilog;
use verilog.vl_types.all;
entity dff_top is
end dff_top;
